-------------------------------------------------------------------------------
-- Declaration
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.fpu_common_p.all;

package fadd_p is

  function fsub (a : fpu_data_t; b : fpu_data_t) return fpu_data_t;
  function fadd (a : fpu_data_t; b : fpu_data_t) return fpu_data_t;

end package;

-------------------------------------------------------------------------------
-- Definition
-------------------------------------------------------------------------------

package body fadd_p is

  function or_nbit (
    a : unsigned;
    n : integer)
    return integer is
  begin
    if unsigned'(a and (shift_left(resize("1", a'length), n) - 1)) = 0 then
      return 0;
    else
      return 1;
    end if;
  end function or_nbit;

  function fadd (
    a : fpu_data_t;
    b : fpu_data_t)
    return fpu_data_t is

    variable fa, fb, fc : float_t;
    variable fbig, fsmall : float_t;

    variable lzc                : integer range 0 to 31;
    variable expdiff            : integer range 0 to 255;
    variable bigfrac, smallfrac : unsigned(23 downto 0);
    variable rawfrac            : unsigned(25 downto 0);

  begin

    fa := float(a);
    fb := float(b);

    ---------------------------------------------------------------------------
    -- sign bit
    ---------------------------------------------------------------------------

    if (fa.sign = "1" and fb.sign = "1")
      or (fa.sign = "1" and (fa.expt & fa.frac) > (fb.expt & fb.frac))
      or (fb.sign = "1" and (fa.expt & fa.frac) < (fb.expt & fb.frac)) then
      fc.sign := "1";
    else
      fc.sign := "0";
    end if;

    ---------------------------------------------------------------------------

    if fa.expt > fb.expt or (fa.expt = fb.expt and fa.frac > fb.frac) then
      fbig   := fa;
      fsmall := fb;
    else
      fbig   := fb;
      fsmall := fa;
    end if;

    expdiff   := to_integer(fbig.expt - fsmall.expt);
    bigfrac   := "1" & fbig.frac & "0";
    if expdiff <= 24 then
      smallfrac := shift_right("1" & fsmall.frac & "0", expdiff)
                   + or_nbit("1" & fsmall.frac & "0", expdiff);
    else
      smallfrac := (others => '0');
    end if;

    if fa.sign /= fb.sign then
      rawfrac := resize(bigfrac, 25) - resize(smallfrac, 25);
    else
      rawfrac :=  resize(smallfrac, 25) + resize(bigfrac, 25);
    end if;

    lzc := leading_zero(rawfrac);

    if lzc = 0 and fbig.expt = 254 then
      fc.expt := (others => '1');
    elsif lzc = 0 then
      fc.expt := fbig.expt + 1;
    elsif lzc = 26 or fbig.expt < lzc then
      fc.expt := (others => '0');
    else
      fc.expt := fbig.expt - (lzc - 1);
    end if;

    if lzc = 0 and fbig.expt = 254 then
      fc.frac := (others => '0');
    elsif lzc = 0 then
      fc.frac := rawfrac(24 downto 2);
    elsif lzc = 26 or fbig.expt < lzc then
      fc.frac := (others => '0');
    else
      fc.frac := shift_left(rawfrac, lzc - 1)(23 downto 1);
    end if;

    ---------------------------------------------------------------------------

    if fa.expt = 0 then
      return b;
    elsif fb.expt = 0 then
      return a;
    elsif fa.expt = 255  and fa.frac /= 0 then
      return VAL_NAN;
    elsif fb.expt = 255 and fb.frac /= 0 then
      return VAL_NAN;
    elsif fa.expt = 255 then
      if fb.expt = 255 and fa.sign /= fb.sign then
        return VAL_NAN;
      else
        return a;
      end if;
    elsif fb.expt = 255 then
      return b;
    else
      return fpu_data(fc);
    end if;

  end function;

  function fsub (
    a : fpu_data_t;
    b : fpu_data_t)
    return fpu_data_t is
    variable nb  : fpu_data_t;
  begin
    nb := (not b(31 downto 31)) & b(30 downto 0);
    return fadd(a, nb);
  end function;
  
end package body fadd_p;
