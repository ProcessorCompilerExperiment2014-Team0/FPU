-------------------------------------------------------------------------------
-- Declaration
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library work;
use work.fpu_common_p.all;

package fsqrt_p is
  component fsqrt is
    port (
      clk: in std_logic;
      a: in std_logic_vector(31 downto 0);
      s: out std_logic_vector(31 downto 0));
  end component;
end package;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

-------------------------------------------------------------------------------
-- Table
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

library work;
use work.fpu_common_p.all;
use work.table_p.all;

entity fsqrt_table_rom is
  port (
    clk: in std_logic;
    en: in std_logic;
    addr: in unsigned(9 downto 0);
    data: out unsigned(35 downto 0));
end fsqrt_table_rom;

architecture behavior of fsqrt_table_rom is

  signal rom: fsqrt_table_t := fsqrt_table;

begin
  process(clk)
  begin
    if rising_edge(clk) then
      if en = '1' then
        data <= ROM(to_integer(addr));
      end if;
    end if;
  end process;
end behavior;

-------------------------------------------------------------------------------
-- Definition
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

library work;
use work.fpu_common_p.all;
use work.fsqrt_p.all;

entity fsqrt is
  port (
    clk: in std_logic;
    a: in std_logic_vector(31 downto 0);
    s: out std_logic_vector(31 downto 0));
end fsqrt;

architecture behavior of fsqrt is
  component fsqrt_table_rom is
    port (
      clk: in std_logic;
      en: in std_logic;
      addr: in unsigned(9 downto 0);
      data: out unsigned(35 downto 0));
  end component;
  signal rom_en: std_logic := '0';
  signal rom_addr: unsigned(9 downto 0);
  signal rom_data: unsigned(35 downto 0);
  type state_t is (NORMAL, CORNER);
  signal state: state_t := CORNER;
  signal state2: state_t := CORNER;
  signal bridge_data: fpu_data_t;
  signal bridge_data2: fpu_data_t;

begin

  table: fsqrt_table_rom port map(
    clk => clk,
    en => rom_en,
    addr => rom_addr,
    data => rom_data);

  fetch: process(clk)
    variable next_state: state_t;
    variable f: float_t;
    variable b: fpu_data_t;
  begin
    if rising_edge(clk) then
      next_state := CORNER;
      if is_metavalue(a) then
        rom_en <= '0';
        b := VAL_NAN;
      else
        f := float(unsigned(a));
        case float_type(f) is
          when NAN =>
            if f.sign = "0" then
              b := VAL_NAN;
            else
              b := VAL_MINUS_NAN;
            end if;
          when INFORMAL =>
            if f.sign = "0" then
              b := VAL_PLUS_ZERO;
            else
              b := VAL_MINUS_ZERO;
            end if;
          when PLUS_INF => b := VAL_PLUS_INF;
          when MINUS_INF => b := VAL_MINUS_NAN;   -- 新たにVAL_MINUS_NANを追加
          when PLUS_ZERO => b := VAL_PLUS_ZERO;
          when MINUS_ZERO => b := VAL_MINUS_ZERO;
          when others =>
            if f.sign = "1" then
              b := VAL_MINUS_NAN;
            else
              next_state := NORMAL;
              rom_en <= '1';
              rom_addr <= (not f.expt(0)) & f.frac(22 downto 14);
              b := unsigned(a);
            end if;
        end case;
      end if;
      bridge_data <= b;
      bridge_data2 <= bridge_data;
      state <= next_state;
      state2 <= state;
    end if;
  end process;

  calc: process(clk)
    variable f, g: float_t;
    variable g_frac_25: unsigned(24 downto 0);
    variable y: unsigned(22 downto 0);
    variable d, n: unsigned(13 downto 0);
    variable ans: unsigned(31 downto 0);
    variable temp_expt: unsigned(7 downto 0);
    variable temp_frac: unsigned(27 downto 0);
  begin
    if rising_edge(clk) then
      case state2 is
        when CORNER =>
          ans := bridge_data2;
        when NORMAL =>
          f := float(bridge_data2);
            g.sign := "0";
            if f.expt >= 127 then
              temp_expt := f.expt - 127;
              temp_expt := shift_right(temp_expt, 1);
              g.expt := 127 + temp_expt;
            else
              temp_expt := 127 - f.expt;
              temp_expt := shift_right(temp_expt+1, 1);
              g.expt := 127 - temp_expt;
            end if;

            y := rom_data(35 downto 13);
            if f.expt(0) = '1' then
              d := '0' & rom_data(12 downto 0);
            else
              d := '1' & rom_data(12 downto 0);
            end if;
            n := f.frac(13 downto 0);
            temp_frac := shift_right(d * n, 14);
            g.frac := y + temp_frac(22 downto 0);
            ans := fpu_data(g);
      end case;
      s <= std_logic_vector(ans);
    end if;
  end process;
end behavior;

            
